module DM(
    input  CLK, RST,
    
)

endmodule